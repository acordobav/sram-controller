class scoreboard;
  int dfifo[$]; // expected data fifo
  int afifo[$]; // address  fifo
  int bfifo[$]; // Burst Length fifo
endclass

`define DUV_PATH top.dut

module whitebox();
  //Define Assertions for WB Interface
  //- Reset
  //- Escritura
  //- Lectura
  //- ...
endmodule
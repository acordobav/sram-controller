interface intf_wb #(parameter dw=32) (input sys_clk, sdram_clk);  //Communicates TB and DUT
	
  //--------------------------------------
  // Wish Bone Interface
  // -------------------------------------      
  logic 				    wb_stb_i;
	logic 				    wb_ack_o;
  logic [25:0] 		  wb_addr_i;
	logic 				    wb_we_i;  // 1 - Write, 0 - Read
	logic [dw-1:0]  	wb_dat_i;
	logic [dw/8-1:0] 	wb_sel_i; // Byte enable
	logic [dw-1:0]  	wb_dat_o;
	logic 				    wb_cyc_i;
  logic [2:0]	 		  wb_cti_i;
  
 	logic sys_clk;
  logic RESETN;

  //--------------------------------------------
  // SDRAM I/F 
  //--------------------------------------------
`ifdef SDR_32BIT
  wire [31:0]      sdr_dq;         // SDRAM Read/Write Data Bus
  wire [3:0]       sdr_dqm ;       // SDRAM DATA Mask
`elsif SDR_16BIT 
  wire [15:0]      sdr_dq;         // SDRAM Read/Write Data Bus
  wire [1:0]       sdr_dqm ;       // SDRAM DATA Mask
`else 
  wire [7:0]       sdr_dq;         // SDRAM Read/Write Data Bus
  wire [0:0]       sdr_dqm;        // SDRAM DATA Mask
`endif

  logic [1:0]       sdr_ba;        // SDRAM Bank Select
  logic [12:0]      sdr_addr;      // SDRAM ADRESS
	logic             sdr_init_done; // SDRAM Init Done 
  
  logic sdram_clk;
  
	logic sdr_cke;
  logic sdr_cs_n;
  logic sdr_ras_n;
  logic sdr_cas_n;
  logic sdr_we_n;

  //--------------------------------------------
  // MODULE PARAMS
  //--------------------------------------------
  logic [1:0]  Req_Depth;
  logic        SDR_Enable;
  logic [12:0] SDR_Mode_Reg;
  logic [3:0]  SDR_tras_d;
  logic [3:0]  SDR_trp_d;
  logic [3:0]  SDR_trcd_d;
  logic [2:0]  SDR_cas;
  logic [3:0]  SDR_trcar_d;
  logic [3:0]  SDR_twr_d;
  logic [11:0] SDR_rf_sh;
  logic [3:0]  SDR_rf_max;

endinterface
